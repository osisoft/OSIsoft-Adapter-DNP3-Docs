<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>OSIsoft Adapter for DNP3 principles of operation </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="OSIsoft Adapter for DNP3 principles of operation ">
    <meta name="generator" content="docfx 2.54.0.0">
    
    <link rel="shortcut icon" href="../../favicon.ico">
    <link rel="stylesheet" href="../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../styles/docfx.css">
    <link rel="stylesheet" href="../../styles/main.css">
    <meta property="docfx:navrel" content="../../toc.html">
    <meta property="docfx:tocrel" content="../toc.html">
    
    <meta property="docfx:rel" content="../../">
    
  </head>
  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              <a class="navbar-brand" href="../../V1/index.html" width="46">
                <img id="logo" src="../../V1/main/V1/images/atlas_icon.png" height="46" width="46" alt="OSIsoft Edge System"> 
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div class="container body-content">
        
        <div id="search-results">
          <div class="search-list"></div>
          <div class="sr-items">
            <p><i class="glyphicon glyphicon-refresh index-loading"></i></p>
          </div>
          <ul id="pagination"></ul>
        </div>
      </div>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="OSIsoftAdapterForDNP3PrinciplesOfOperation">
<h1 id="osisoft-adapter-for-dnp3-principles-of-operation" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="5" sourceendlinenumber="5">OSIsoft Adapter for DNP3 principles of operation</h1>

<h2 id="connectivity-and-interoperability" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="7" sourceendlinenumber="7">Connectivity and Interoperability</h2>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="8" sourceendlinenumber="8">The DNP3 Adapter may connect to one or more DNP3 compliant outstations via TCP/IP connections. The total number of outstations that the DNP3 Adapter may connect to will vary across different installation environments.  </p>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="10" sourceendlinenumber="13">The DNP3 Adapter is designed to operate with Level 1 (DNP3–L1) compliance, which defines minimum requirements for all DNP3 compliant devices. 
However, the adapter does make use of some Level 2, Level 3, and Level 4 functions. Some DNP3 compliant devices may not support these same features.<br>Any functionality described in this documentation that is not required for Level 1 compliance will be noted as such. 
Please check the outstation documentation prior to using these features, as the adapter will need to be configured to only use the supported features of the outstation.  </p>
<h2 id="adapter-configuration" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="15" sourceendlinenumber="15">Adapter Configuration</h2>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="17" sourceendlinenumber="17">In order for the DNP3 Adapter to start data collection, you need to configure the adapter by defining the following:</p>
<ul sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="19" sourceendlinenumber="21">
<li sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="19" sourceendlinenumber="19">Data source: Provide the information required to connect to your DNP3 compliant outstations. </li>
<li sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="20" sourceendlinenumber="20">Data selection: Select the DNP points on the outstations you want the adapter to collect data from.</li>
<li sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="21" sourceendlinenumber="21">Logging: Set up the logging attributes to manage the adapter logging behavior.</li>
</ul>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="23" sourceendlinenumber="23">For more infomation, see <a class="xref" href="../Configuration/OSIsoft%20Adapter%20for%20DNP3%20data%20source%20configuration.html" data-raw-source="[OSIsoft Adapter for DNP3 data source configuration](xref:OSIsoftAdapterForDNP3DataSourceConfiguration)" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="23" sourceendlinenumber="23">OSIsoft Adapter for DNP3 data source configuration</a> and <a class="xref" href="../Configuration/OSIsoft%20Adapter%20for%20DNP3%20data%20selection%20configuration.html" data-raw-source="[OSIsoft Adapter for DNP3 data selection configuration](xref:OSIsoftAdapterForDNP3DataSelectionConfiguration)" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="23" sourceendlinenumber="23">OSIsoft Adapter for DNP3 data selection configuration</a>.</p>
<h2 id="stream-creation" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="25" sourceendlinenumber="25">Stream creation</h2>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="26" sourceendlinenumber="26">The DNP3 adapter creates types at startup. One stream is created for every selected DNP point represented by an item in the data selection configuration. Each stream contains two properties:</p>
<table sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="28" sourceendlinenumber="31">
<thead>
<tr>
<th>Property name</th>
<th>Data type</th>
<th>Description</th>
</tr>
</thead>
<tbody>
<tr>
<td>Timestamp</td>
<td>DateTime</td>
<td>Timestamp of the value update for the DNP point.</td>
</tr>
<tr>
<td>Value</td>
<td>Depenent on the data selection configuration</td>
<td>Value of the DNP point</td>
</tr>
</tbody>
</table>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="33" sourceendlinenumber="34">Each stream will have a unique identifier, called a Stream ID, which can be specified by the user in the data selection configuration. 
If the Stream ID is not specified, the adapter will use the DefaultStreamIdPattern in the data source configuration to determine the Stream ID. </p>
<h3 id="discovery" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="36" sourceendlinenumber="36">Discovery</h3>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="37" sourceendlinenumber="41">The DNP3 adapter can discover points on your DNP3 outstation by performing an <a href="#Integrity-scan" data-raw-source="[*integrity scan*](#Integrity-scan)" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="37" sourceendlinenumber="37"><em>integrity scan</em></a>. 
Discovery will populate your data selection configuration with items that represent points on the outstation. 
These items will default as unselected, so the user may make changes to these items before selecting them. 
The adapter can only discover points that are assigned to Class 0, Class 1, Class 2, or Class 3 on the outstation.
Discovery may be expensive in terms of bandwidth and outstation resources, so the adapter will only perform discovery for an outstation when the following criteria is met: </p>
<ul sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="43" sourceendlinenumber="45">
<li sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="43" sourceendlinenumber="43">The outstation is configured in the data source configuration.</li>
<li sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="44" sourceendlinenumber="44">The adapter is configured to perform an integrity scan for that outstation. </li>
<li sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="45" sourceendlinenumber="45">The data selection configuration contains no items that correlate to that outstation, selected or unselected.</li>
</ul>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="47" sourceendlinenumber="51">To discover a new outstation, simply add the outstation to the data source configuration and configure an integrity scan to run periodically or on startup. 
The adapter will use the first integrity scan as a means for discovery. 
To configure a new outstation without triggering a discovery, you can add one or more selection items to correspond with the outstation. 
The items may be selected or unselected. 
Alternatively, you can configure the outstation behavior so that no integrity scan will be performed. Without an integrity scan, discovery will not be possible. </p>
<h2 id="data-collection" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="53" sourceendlinenumber="53">Data collection</h2>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="54" sourceendlinenumber="54">The DNP3 adapter can collect two different types of data from DNP3 compliant outstations: <em>static</em> data and <em>event</em> data.</p>
<h3 id="static-data" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="56" sourceendlinenumber="56">Static data</h3>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="57" sourceendlinenumber="62">The DNP3 specification defines static data as the current value of a DNP point at the time of a request. 
The DNP3 adapter may be configured to request static data by polling the outstation(s) for a range of points that share an object group and variation,
 which are configured in the data selection configuration. 
Static data will be reported with the current time of the adapter machine. 
When polling for static data at predefined rate, it is possible that quickly changing data may be missed by the adapter. 
It is also possible that the adapter will receive multiple values representing the same event but with different timestamps. </p>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="64" sourceendlinenumber="69">The adapter makes a request for the current value of specific points as configured in the Data Selection configuration file. 
The adapter will request this data via a range scan, which will request the static data for a range of point indices that share a group and variation,
 as configured in the data selection configuration.
The outstation should report the current value of each point, but the outstation is not required to report using the requested object variation. 
If the outstation responds with a different variation than what the adapter has requested, the adapter will still send the data it receives.
This could lead to differences in the reported value versus what is expected in terms of precision and status. </p>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="71" sourceendlinenumber="73">Support for requesting static data for DNP3 points via a range scan is at least a Level 2 function, and some groups and variations may be considered L3 or L4 functionality.
Because of this, it is important to verify that your outstation supports this functionality before configuring the adapter to collect data in this manner. 
Some DNP3-L1 compliant outstations may optionally support this type of scan. </p>
<h3 id="event-data" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="75" sourceendlinenumber="75">Event data</h3>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="76" sourceendlinenumber="85">The DNP3 specification defines event data as the information that is retained regarding an event. 
An event is defined by the DNP3 specification as the occurrence of something significant happening. 
What constitutes an event may vary depending on the implementation of the outstation. 
Typically, an event will result in a value change for a DNP point,
 although it is possible for an event to occur that does not change the value of any point on the outstation. 
Event data is saved at the outstation(s) and should be kept until the adapter confirms that it has received the event object.<br>The event object is the description of the event that the adapter should receive from the outstation(s). 
The event object may contain the value, time, and status code relating to the event and corresponding point. 
The exact information contained in the object will be dependent on both the point type and variation,
 which are defined in the DNP3 specification.  </p>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="87" sourceendlinenumber="89">DNP3 events belong to one of three different classes of data: <em>Class 1</em>, <em>Class 2</em>, or <em>Class 3</em>. 
These event classes may be used to group events by priority,
 though neither the DNP3 adapter nor the DNP3 specification assign significance to the three event classes. </p>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="91" sourceendlinenumber="91">According to the DNP3 specification, all DNP3 – L1 compliant outstations shall accept read requests for event class data.  </p>
<h4 id="event-scans" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="93" sourceendlinenumber="93">Event Scans</h4>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="94" sourceendlinenumber="96">The adapter may be configured to request event data via an <em>event scan</em>. 
During an <em>event scan</em>, the adapter will poll the outstation(s) for the event data from each of the configured event classes. 
The event classes and the polling interval may be configured in the <a class="xref" href="../Configuration/OSIsoft%20Adapter%20for%20DNP3%20data%20source%20configuration.html#OutstationBehavior-Parameters" data-raw-source="[data source configuration](xref:OSIsoftAdapterForDNP3DataSourceConfiguration#OutstationBehavior-Parameters)" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="96" sourceendlinenumber="96">data source configuration</a>.</p>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="98" sourceendlinenumber="105"><em>Event scans</em> offer several advantages over polling for static data. 
When polling for static data, it is possible to miss value changes for points on the outstation;
 however, <em>event scans</em> will ensure that each outstation reports every event to the adapter. 
Similarly, even when polling quickly, some events could be missed if they do not change the value of the DNP point. 
If bandwidth is a concern, the adapter may make efficient use of the network by only requesting event data. 
When polling for static data, the outstation may report unchanging data unnecessarily, whereas <em>event scans</em> should only return new events. 
It is important to configure the adapter to perform Event Scans at an interval that is not long enough to allow the outstations’ event buffers to become full. 
Refer to the documentation for each specific outstation to determine what constitutes an event and how much time it will take before the buffer becomes full. </p>
<h4 id="unsolicited-events" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="107" sourceendlinenumber="107">Unsolicited Events</h4>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="108" sourceendlinenumber="109">In addition to the <em>event scans</em> above, the adapter may be configured to receive <em>unsolicited</em> responses containing event data. 
An unsolicited response is a message sent from an outstation that the adapter did not explicitly request. </p>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="111" sourceendlinenumber="113">If the adapter is configured to receive unsolicited data, outstations that support sending unsolicited data should report event data to the adapter as it occurs. 
This could eliminate the need for the adapter to poll the outstation(s) for data. 
The decision to configure the adapter to receive unsolicited data, or to perform Event Scans should be carefully considered.  </p>
<h3 id="integrity-scans" sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="115" sourceendlinenumber="115">Integrity Scans</h3>
<p sourcefile="V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md" sourcestartlinenumber="116" sourceendlinenumber="123">The DNP3 adapter can be configured to perform an <em>integrity scan</em> on startup,
 when the outstation&#39;s event buffer overflows, and/or at a defined interval.
During an <em>integrity scan</em>, the adapter will poll the outstation(s) for events,
 then the current value of all points that are assigned to one of the event classes (or class 0).
The adapter performs an integrity scan by polling Object Group 60.
If bandwidth or outstation performance is a concern, carefully consider the value of an integrity scan, as the outstation may respond with data for many more points than the adapter is configured to collect data for. 
The adapter will simply discard any data that it receives without a corresponding data selection item. 
To retrieve the current value of any points not assigned to an event class, the adapter will need to perform a <em>static scan</em>.</p>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                  <li>
                    <a href="https://github.com/osisoft/OSIsoft-Adapter-DNP3-Docs/blob/master/V1/OSIsoft Adapter for DNP3 overview/OSIsoft Adapter for DNP3 principles of operation.md/#L1" class="contribution-link">Improve this Doc</a>
                  </li>
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
              <!-- <p><a class="back-to-top" href="#top">Back to top</a><p> -->
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>© 2020 - OSIsoft, LLC.</span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../styles/main.js"></script>
  </body>
</html>
